package constants is

    -- Lattice iCEStick40 clock frequency
    constant clock_frequency : real := 12.0e6;

    -- how long each LED should be lit in milliseconds
    constant led_pulse_time_ms : natural := 250;

end package;